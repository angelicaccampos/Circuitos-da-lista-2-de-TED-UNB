CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
210 120 30 250 10
190 80 1286 747
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
358 176 471 273
9437202 0
0
6 Title:
5 Name:
0
0
0
10
13 Logic Switch~
5 307 322 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3536 0 0
2
45229.7 0
0
13 Logic Switch~
5 305 276 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4597 0 0
2
45229.7 0
0
13 Logic Switch~
5 303 223 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3835 0 0
2
45229.7 0
0
13 Logic Switch~
5 302 172 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3670 0 0
2
45229.7 0
0
14 Logic Display~
6 494 214 0 1 2
29 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5616 0 0
2
45229.7 0
0
8 2-In OR~
219 449 232 0 3 22
0 4 7 6
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U2A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
9323 0 0
2
45229.7 0
0
12 2-In NOR:DM~
219 463 181 0 3 22
0 5 2 9
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
317 0 0
2
45229.7 0
0
5 7415~
219 404 267 0 4 22
0 2 5 8 7
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 1 0
1 U
3108 0 0
2
45229.7 0
0
5 7415~
219 403 223 0 4 22
0 5 2 3 4
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 1 0
1 U
4299 0 0
2
45229.7 0
0
14 Logic Display~
6 494 162 0 1 2
46 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9672 0 0
2
45229.7 0
0
12
1 0 2 0 0 4096 0 8 0 0 2 4
380 258
333 258
333 222
334 222
0 2 2 0 0 8336 0 0 7 3 0 3
334 223
334 190
433 190
1 2 2 0 0 0 0 3 9 0 0 2
315 223
379 223
3 1 3 0 0 8320 0 9 1 0 0 4
379 232
361 232
361 322
319 322
4 1 4 0 0 4224 0 9 6 0 0 2
424 223
436 223
0 2 5 0 0 4224 0 0 8 12 0 3
320 172
320 267
380 267
3 1 6 0 0 4224 0 6 5 0 0 2
482 232
494 232
4 2 7 0 0 8320 0 8 6 0 0 3
425 267
436 267
436 241
1 3 8 0 0 4224 0 2 8 0 0 2
317 276
380 276
3 1 9 0 0 4224 0 7 10 0 0 3
484 181
494 181
494 180
0 1 5 0 0 0 0 0 7 12 0 2
379 172
433 172
1 1 5 0 0 0 0 4 9 0 0 3
314 172
379 172
379 214
6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
502 206 519 230
506 209 514 225
1 G
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
503 154 520 178
507 157 515 173
1 R
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
271 263 288 287
275 266 283 282
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
272 309 289 333
276 312 284 328
1 D
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
269 211 286 235
273 214 281 230
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
270 160 287 184
274 163 282 179
1 A
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
