CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
270 80 30 250 10
176 80 1286 747
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
12
13 Logic Switch~
5 319 281 0 1 11
0 2
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
45229.6 0
0
13 Logic Switch~
5 319 237 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
45229.6 0
0
13 Logic Switch~
5 319 196 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3124 0 0
2
45229.6 0
0
13 Logic Switch~
5 320 156 0 1 11
0 12
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3421 0 0
2
45229.6 0
0
9 2-In AND~
219 516 233 0 3 22
0 6 4 5
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
8157 0 0
2
45229.6 0
0
8 2-In OR~
219 559 242 0 3 22
0 5 2 7
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
5572 0 0
2
45229.6 0
0
9 Inverter~
13 463 242 0 2 22
0 2 4
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
8901 0 0
2
45229.6 0
0
8 2-In OR~
219 459 196 0 3 22
0 3 8 6
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
7361 0 0
2
45229.6 0
0
9 2-In AND~
219 417 205 0 3 22
0 10 9 8
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
4747 0 0
2
45229.6 0
0
9 2-In AND~
219 617 164 0 3 22
0 12 7 11
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
972 0 0
2
45229.6 0
0
14 Logic Display~
6 653 144 0 1 2
12 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3472 0 0
2
45229.6 0
0
9 Inverter~
13 365 196 0 2 22
0 3 10
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
9998 0 0
2
45229.6 0
0
13
3 2 0 0 0 0 0 9 8 0 0 2
438 205
446 205
1 1 2 0 0 12432 0 7 1 0 0 4
448 242
447 242
447 281
331 281
1 0 3 0 0 8320 0 8 0 0 11 4
446 187
446 171
344 171
344 196
2 2 4 0 0 4224 0 7 5 0 0 2
484 242
492 242
3 1 5 0 0 4224 0 5 6 0 0 2
537 233
546 233
3 1 6 0 0 4224 0 8 5 0 0 2
492 196
492 224
3 2 7 0 0 4224 0 6 10 0 0 3
592 242
592 173
593 173
0 2 2 0 0 4224 0 0 6 2 0 4
447 280
543 280
543 251
546 251
1 2 9 0 0 4224 0 2 9 0 0 3
331 237
393 237
393 214
2 1 10 0 0 12416 0 12 9 0 0 4
386 196
378 196
378 196
393 196
1 1 3 0 0 0 0 3 12 0 0 2
331 196
350 196
3 1 11 0 0 4224 0 10 11 0 0 3
638 164
653 164
653 162
1 1 12 0 0 4224 0 4 10 0 0 4
332 156
578 156
578 155
593 155
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
659 134 688 158
669 142 677 158
1 S
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
271 261 300 285
281 269 289 285
1 D
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
272 218 301 242
282 226 290 242
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
272 176 301 200
282 184 290 200
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
272 135 301 159
282 143 290 159
1 A
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
