CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
30 160 30 260 10
158 80 1286 747
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
326 176 439 273
9437202 0
0
6 Title:
5 Name:
0
0
0
12
13 Logic Switch~
5 68 385 0 1 11
0 4
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V

%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8396 0 0
2
45227.3 0
0
13 Logic Switch~
5 70 294 0 1 11
0 2
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V

%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3685 0 0
2
45227.3 0
0
13 Logic Switch~
5 70 195 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V

%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7849 0 0
2
45227.3 0
0
8 4-In OR~
219 338 298 0 5 22
0 12 10 9 8 11
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U3A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 3 0
1 U
6343 0 0
2
45227.3 0
0
14 Logic Display~
6 384 260 0 1 2
24 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7376 0 0
2
45227.3 0
0
9 Inverter~
13 166 340 0 2 22
0 4 5
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 4 0
1 U
9156 0 0
2
45227.3 0
0
9 Inverter~
13 167 252 0 2 22
0 2 6
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 4 0
1 U
5776 0 0
2
45227.3 0
0
9 Inverter~
13 159 195 0 2 22
0 3 7
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
7207 0 0
2
45227.3 0
0
5 7415~
219 268 394 0 4 22
0 4 2 3 8
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 2 0
1 U
4459 0 0
2
45227.3 0
0
5 7415~
219 268 349 0 4 22
0 5 6 3 9
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 1 0
1 U
3760 0 0
2
45227.3 0
0
5 7415~
219 269 294 0 4 22
0 7 2 5 10
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 1 0
1 U
754 0 0
2
45227.3 0
0
5 7415~
219 270 204 0 4 22
0 7 4 6 12
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 1 0
1 U
9767 0 0
2
45227.3 0
0
19
0 2 2 0 0 4096 0 0 9 9 0 3
144 294
144 394
244 394
3 0 3 0 0 4096 0 9 0 0 4 4
244 403
95 403
95 358
96 358
0 1 4 0 0 4096 0 0 9 11 0 2
151 385
244 385
0 3 3 0 0 4224 0 0 10 14 0 3
96 195
96 358
244 358
2 3 5 0 0 4224 0 6 11 0 0 4
187 340
243 340
243 303
245 303
0 2 4 0 0 4224 0 0 12 11 0 4
120 385
120 208
246 208
246 204
0 3 6 0 0 8192 0 0 12 8 0 3
191 252
191 213
246 213
2 2 6 0 0 8320 0 7 10 0 0 4
188 252
191 252
191 349
244 349
0 2 2 0 0 4224 0 0 11 12 0 2
144 294
245 294
0 1 7 0 0 4224 0 0 11 13 0 3
221 195
221 285
245 285
1 1 4 0 0 0 0 1 6 0 0 3
80 385
151 385
151 340
1 1 2 0 0 0 0 2 7 0 0 4
82 294
144 294
144 252
152 252
2 1 7 0 0 0 0 8 12 0 0 2
180 195
246 195
1 1 3 0 0 0 0 3 8 0 0 2
82 195
144 195
4 4 8 0 0 8320 0 9 4 0 0 4
289 394
314 394
314 312
321 312
4 3 9 0 0 8320 0 10 4 0 0 4
289 349
302 349
302 303
321 303
4 2 10 0 0 4224 0 11 4 0 0 2
290 294
321 294
5 1 11 0 0 8320 0 4 5 0 0 3
371 298
384 298
384 278
4 1 12 0 0 8320 0 12 4 0 0 4
291 204
300 204
300 285
321 285
4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
388 248 413 272
396 256 404 272
1 S
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
33 367 62 391
43 375 51 391
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
32 282 61 306
42 290 50 306
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
34 175 63 199
44 183 52 199
1 A
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 1e-06 1e-07 1e-07
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
