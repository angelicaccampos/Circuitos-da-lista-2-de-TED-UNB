CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
220 120 30 370 10
146 80 1286 747
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
314 176 427 273
9437202 0
0
6 Title:
5 Name:
0
0
0
10
13 Logic Switch~
5 260 277 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V

%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5283 0 0
2
45227.3 0
0
13 Logic Switch~
5 259 214 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V

%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6874 0 0
2
45227.3 0
0
13 Logic Switch~
5 260 177 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V

%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5305 0 0
2
45227.3 1
0
5 4073~
219 359 264 0 4 22
0 2 6 5 3
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 4 0
1 U
34 0 0
2
45227.3 0
0
9 Inverter~
13 307 264 0 2 22
0 4 6
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
969 0 0
2
45227.3 0
0
9 Inverter~
13 305 196 0 2 22
0 7 2
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
8402 0 0
2
45227.3 0
0
14 Logic Display~
6 401 230 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3751 0 0
2
5.90097e-315 0
0
14 Logic Display~
6 400 187 0 1 2
23 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4292 0 0
2
45227.3 2
0
14 Logic Display~
6 400 146 0 1 2
11 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6118 0 0
2
45227.3 3
0
9 2-In AND~
219 359 205 0 3 22
0 2 4 8
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
34 0 0
2
45227.3 4
0
10
0 1 2 0 0 4224 0 0 4 7 0 3
329 196
329 255
335 255
4 1 3 0 0 4224 0 4 7 0 0 3
380 264
401 264
401 248
1 0 4 0 0 8192 0 5 0 0 6 3
292 264
281 264
281 214
1 3 5 0 0 4224 0 1 4 0 0 3
272 277
335 277
335 273
2 2 6 0 0 4224 0 5 4 0 0 2
328 264
335 264
1 2 4 0 0 4224 0 2 10 0 0 2
271 214
335 214
2 1 2 0 0 0 0 6 10 0 0 2
326 196
335 196
0 1 7 0 0 4096 0 0 6 9 0 3
282 177
282 196
290 196
1 1 7 0 0 12432 0 3 9 0 0 4
272 177
282 177
282 164
400 164
3 1 8 0 0 4224 0 10 8 0 0 2
380 205
400 205
6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
232 264 249 287
236 268 244 283
1 R
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
226 200 249 223
229 204 245 219
2 TF
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
225 163 250 186
229 167 245 182
2 TD
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
411 226 434 250
414 228 430 244
2 Sc
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
411 182 434 206
414 184 430 200
2 Sb
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
409 141 432 165
412 143 428 159
2 Sa
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
