CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
60 120 30 180 10
127 80 1286 747
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
295 176 408 273
9437202 0
0
6 Title:
5 Name:
0
0
0
14
13 Logic Switch~
5 154 206 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9592 0 0
2
45227.3 0
0
13 Logic Switch~
5 157 291 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8748 0 0
2
5.90097e-315 0
0
14 Logic Display~
6 386 367 0 1 2
12 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7168 0 0
2
45227.3 0
0
9 Inverter~
13 236 413 0 2 22
0 5 4
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 3 0
1 U
631 0 0
2
45227.3 0
0
9 Inverter~
13 236 371 0 2 22
0 3 9
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 3 0
1 U
9466 0 0
2
45227.3 0
0
9 Inverter~
13 236 337 0 2 22
0 5 8
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
3266 0 0
2
45227.3 0
0
5 4071~
219 345 389 0 3 22
0 7 2 6
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U2B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
7693 0 0
2
45227.3 0
0
5 4081~
219 302 421 0 3 22
0 4 3 2
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U1D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 1 0
1 U
3723 0 0
2
45227.3 0
0
5 4081~
219 301 362 0 3 22
0 8 9 7
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 1 0
1 U
3440 0 0
2
45227.3 0
0
14 Logic Display~
6 385 221 0 1 2
21 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6263 0 0
2
45227.3 0
0
9 Inverter~
13 235 224 0 2 22
0 3 13
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
4900 0 0
2
45227.3 0
0
5 4071~
219 343 245 0 3 22
0 12 11 10
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U2A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
8783 0 0
2
45227.3 0
0
5 4081~
219 302 282 0 3 22
0 5 3 11
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 1 0
1 U
3221 0 0
2
45227.3 0
0
5 4081~
219 301 215 0 3 22
0 5 13 12
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
3215 0 0
2
45227.3 0
0
18
3 2 2 0 0 4224 0 8 7 0 0 3
323 421
323 398
332 398
0 2 3 0 0 4224 0 0 8 18 0 3
179 291
179 430
278 430
2 1 4 0 0 8320 0 4 8 0 0 3
257 413
257 412
278 412
0 1 5 0 0 4224 0 0 4 16 0 3
188 206
188 413
221 413
3 1 6 0 0 4224 0 7 3 0 0 3
378 389
386 389
386 385
3 1 7 0 0 4224 0 9 7 0 0 3
322 362
322 380
332 380
2 1 8 0 0 8320 0 6 9 0 0 3
257 337
257 353
277 353
2 2 9 0 0 4224 0 5 9 0 0 2
257 371
277 371
0 1 3 0 0 0 0 0 5 18 0 3
210 291
210 371
221 371
0 1 5 0 0 16 0 0 6 16 0 3
198 206
198 337
221 337
3 1 10 0 0 4224 0 12 10 0 0 3
376 245
385 245
385 239
3 2 11 0 0 4224 0 13 12 0 0 3
323 282
323 254
330 254
3 1 12 0 0 4224 0 14 12 0 0 3
322 215
322 236
330 236
0 2 3 0 0 0 0 0 13 18 0 2
219 291
278 291
0 1 5 0 0 0 0 0 13 16 0 3
268 206
268 273
278 273
1 1 5 0 0 128 0 1 14 0 0 2
166 206
277 206
2 2 13 0 0 4224 0 11 14 0 0 2
256 224
277 224
1 1 3 0 0 128 0 2 11 0 0 3
169 291
220 291
220 224
4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
398 359 425 383
404 363 418 379
2 R1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
397 212 424 236
403 217 417 233
2 R2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
125 279 143 303
130 284 137 300
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
123 198 141 222
128 203 135 219
1 A
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
