CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
70 140 30 340 10
168 80 1286 747
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
336 176 449 273
9437202 0
0
6 Title:
5 Name:
0
0
0
10
13 Logic Switch~
5 104 267 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9172 0 0
2
5.90097e-315 0
0
13 Logic Switch~
5 102 210 0 1 11
0 2
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7100 0 0
2
5.90097e-315 0
0
13 Logic Switch~
5 102 173 0 1 11
0 6
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3820 0 0
2
5.90097e-315 0
0
14 Logic Display~
6 362 216 0 1 2
31 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7678 0 0
2
5.90097e-315 0
0
9 Inverter~
13 182 267 0 2 22
0 8 7
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 3 0
1 U
961 0 0
2
5.90097e-315 0
0
9 Inverter~
13 222 210 0 2 22
0 2 9
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
3178 0 0
2
5.90097e-315 0
0
9 Inverter~
13 220 173 0 2 22
0 6 10
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
3409 0 0
2
5.90097e-315 0
0
8 2-In OR~
219 324 242 0 3 22
0 5 4 3
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U2A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3951 0 0
2
5.90097e-315 0
0
5 7415~
219 280 279 0 4 22
0 7 6 2 4
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 1 0
1 U
8885 0 0
2
5.90097e-315 0
0
5 7415~
219 281 210 0 4 22
0 10 9 8 5
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 1 0
1 U
3780 0 0
2
5.90097e-315 0
0
12
0 3 2 0 0 8320 0 0 9 11 0 3
130 210
130 288
256 288
3 1 3 0 0 8336 0 8 4 0 0 3
357 242
362 242
362 234
4 2 4 0 0 4224 0 9 8 0 0 3
301 279
301 251
311 251
4 1 5 0 0 4224 0 10 8 0 0 3
302 210
302 233
311 233
0 2 6 0 0 8320 0 0 9 12 0 3
146 173
146 279
256 279
2 1 7 0 0 4224 0 5 9 0 0 4
203 267
243 267
243 270
256 270
0 3 8 0 0 8320 0 0 10 10 0 4
157 267
157 223
257 223
257 219
2 2 9 0 0 12416 0 6 10 0 0 4
243 210
242 210
242 210
257 210
2 1 10 0 0 8320 0 7 10 0 0 4
241 173
247 173
247 201
257 201
1 1 8 0 0 0 0 1 5 0 0 2
116 267
167 267
1 1 2 0 0 0 0 2 6 0 0 2
114 210
207 210
1 1 6 0 0 0 0 3 7 0 0 2
114 173
205 173
4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
370 190 385 214
373 192 381 208
1 S
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
74 254 89 278
77 256 85 272
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
73 202 88 226
76 204 84 220
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
73 160 88 184
76 162 84 178
1 A
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
